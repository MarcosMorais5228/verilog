module NOT (input A, output F);
    nand(F,A,A)
    
endmodule